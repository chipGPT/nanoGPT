
// macros
// bit width
`define EXP_SIZE    4
`define MNT_SIZE    3   
`define DATA_SIZE   8
`define ADDR_SIZE   20
// input config
`define INPUT_NUM   12
`define ROW_NUM     24
// address
`define ADDR_BASE   0
`define ADDR_OFFU   1'b1

