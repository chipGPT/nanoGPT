// Copyright (c) 2024, Saligane's Group at University of Michigan and Google Research
//
// Licensed under the Apache License, Version 2.0 (the "License");

// you may not use this file except in compliance with the License.

// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// macros
// bit width
`define EXP_SIZE    4
`define MNT_SIZE    3   
`define DATA_SIZE   8
`define ADDR_SIZE   20
// input config
`define INPUT_NUM   12
`define ROW_NUM     24
// address
`define ADDR_BASE   0
`define ADDR_OFFU   1'b1

